module PC();
	input clk;
	input [31:0] prox_endereco